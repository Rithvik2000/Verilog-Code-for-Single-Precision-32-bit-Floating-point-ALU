`timescale 1ns / 100ps


module TB_for_ALU #(parameter N = 32)();
reg [N-1:0] A;
reg [N-1:0] B;
reg [2:0] Select;

wire [N-1:0] OUT;
wire Underflow,Overflow;

FP_ALU a1(A,B,Select,OUT,Underflow,Overflow);





initial begin

//$monitor(" a = %f | b = %f| pp = %f| CLK = %B |RST = %b|acc = %f |Un = %b |Ov = %b",
// A,B,Partial_Product,CLK,RST,ACC,Underflow,Overflow);
 #5
Select = 1;

#30

A =32'b11000000011000111100000000000000 ; 
B =32'b01000000101101000000000000000000 ;

#30

A =32'b00111111100111000000000000000000 ; 
B =32'b11111110101000000000000000000000 ;

#30


A =32'b01010101010101010101110101010101;
B =32'b01010101010101010101110101010101;

#30

A =32'b01000001010101011101010101010101;
B =32'b01000100110101010101010101010101;

#30

A =32'b01000001011111010101010101010101;
B =32'b01000011110101010101010101010101;

#30

A =32'b00000001100000000000000000000000;
B =32'b00000001100000000000000000000000;

#30

A =32'b11111111011111111111111111111111;
B =32'b11111111011111111111111111111111;

#30


Select = 2;

#30

A =32'b11000000011000111100000000000000 ; 
B =32'b01000000101101000000000000000000 ;

#30

A =32'b00111111100111000000000000000000 ; 
B =32'b11111110101000000000000000000000 ;




#30


A =32'b01000000010111010101110101010101;
B =32'b01000000011101010101110101010101;

#30

A =32'b01000000010101011101010101010101;
B =32'b01000000010101010101010101010101;

#30

A =32'b01010101011111010101010101010101;
B =32'b01010111110101010101010101010101;



Select = 3;
#30

A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b01000011011111100000000001111111;
B =32'b11000011011111111000000001111111;
#40

#30
A =32'b0100101011111111111111111010101;
B =32'b0011101010101010101110101010101;

#30


A =32'b01000111010101011101010101010101;
B =32'b01000101100000000101010101010101;

#30

A =32'b00000000000000000000000000000000;
B =32'b01000101100000000101010101010101;

#30


A =32'b11111111111111111111111111111111;
B =32'b11111111111111111111111111111111;

#30


A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b01000011011111100000000001111111;
B =32'b11000011011111111000000001111111;



#30
A =32'b01000101011111111111111111010101;
B =32'b11010101010101010101110101010101;

#30
A =32'b00000000000001000000000000000000;
B =32'b10000000000000010000000000000000;

#30
A =32'b01000101010101011101010101010101;
B =32'b11000000000000000101010101010101;

#30
A =32'b01010101011111111111111111010101;
B =32'b01010101010101010101110101010101;

#30
A =32'b01010101010101011101010101010101;
B =32'b01010101100000000101010101010101;


Select = 4;
#30

A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b01000011011111100000000001111111;
B =32'b11000011011111111000000001111111;
#40

#30
A =32'b0100101011111111111111111010101;
B =32'b0011101010101010101110101010101;

#30


A =32'b01000111010101011101010101010101;
B =32'b01000101100000000101010101010101;

#30

A =32'b00000000000000000000000000000000;
B =32'b01000101100000000101010101010101;

#30


A =32'b01000111101110000000000000000000;
B =32'b11000111101101000000000000000000;

#30


A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b01000011011111100000000001111111;
B =32'b11000011011111111000000001111111;



#30
A =32'b01000101011111111111111111010101;
B =32'b11010101010101010101110101010101;

#30
A =32'b00000000000001000000000000000000;
B =32'b10000000000000010000000000000000;

#30
A =32'b01000101010101011101010101010101;
B =32'b11000000000000000101010101010101;

#30
A =32'b01010101011111111111111111010101;
B =32'b01010101010101010101110101010101;

#30
A =32'b01010101010101011101010101010101;
B =32'b01010101100000000101010101010101;



Select = 5;
#30

A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b01000011011111100000000001111111;
B =32'b11000011011111111000000001111111;
#40

#30
A =32'b0100101011111111111111111010101;
B =32'b0011101010101010101110101010101;

#30


A =32'b01000111010101011101010101010101;
B =32'b01000101100000000101010101010101;

#30

A =32'b00000000000000000000000000000000;
B =32'b01000101100000000101010101010101;

#30


A =32'b01000111101110000000000000000000;
B =32'b11000111101101000000000000000000;

#30


A =32'b11000101100001111111100000000000;
B =32'b01000001100000000000001111100000;

#30


A =32'b11000011011111111000000001111111;
B =32'b11000011011111111000000001111111;



#30
A =32'b01000101011111111111111111010101;
B =32'b11010101010101010101110101010101;

#30
A =32'b00000000000001000000000000000000;
B =32'b10000000000000010000000000000000;

#30
A =32'b01000101010101011101010101010101;
B =32'b11000000000000000101010101010101;

#30
A =32'b01010101010101010101110101010101;
B =32'b01010101010101010101110101010101;

#30
A =32'b01010101010101011101010101010101;
B =32'b01010101100000000101010101010101;

#30


$finish;
end

endmodule
